module SignExt(BusImm, Imm26, Ctrl); 
   output [63:0] BusImm; 
   input [25:0]  Imm26; 
   input [2:0]	 Ctrl; 
   
   reg [63:0] BusImm;
   always @(*)
      begin
	case (Ctrl)
	3'b000: BusImm = {{52{1'b0}}, Imm26[21:10]}; //I-type: 12 bit immedite (zero extend)
	3'b001: BusImm = {{55{Imm26[20]}}, Imm26[20:12]};  //D-type: 9 bit address
	3'b010: BusImm = {{38{Imm26[25]}}, Imm26}; //B-type: 26 bit address
	3'b011: BusImm = {{45{Imm26[23]}}, Imm26[23:5]}; //CB-type: 19 bit address
	default: BusImm = {{46{1'b0}}, Imm26[22:5]};   //default is movz
	endcase
      end
   
endmodule
